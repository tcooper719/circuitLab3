module halfAdder (output S, C, input x, y);
    xor (S, x, y);
    and (C, x, y);
endmodule